module inverter (inp, op);

input inp; 
output op;

assign op = ~inp; 

endmodule
