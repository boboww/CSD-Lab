module Lab5_Cont(
    );


endmodule
