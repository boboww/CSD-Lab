module Lab5_Cont(
    );

//So this would be where we would have the sequntial code (states)
//if they needed to go here. 

//I currently have the sequential stuff in the main Lab5.v file and
//it would probably be simpler to keep everything there if possible. 

//Might be messier though.

//Move stuff here if neccessary. Just look at the "other group's"
//for inspiration 

endmodule
